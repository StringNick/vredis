module vredis


pub fn should_retry(err IError, retry_timeout bool) bool {
	if err == nil_value {
		return false
	}

	return false
}
