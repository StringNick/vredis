module vredis

fn test_q() {
	//new_client()
	mut cl := new_client(Options{})
	eprintln('client $cl')
}
