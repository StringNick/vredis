module pool


fn test_q() {}
